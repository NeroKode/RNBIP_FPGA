`timescale 1ns / 1ps

module MemCache(
    input [7:0] Address,
               //inout [7:0] DataBus,
                input [7:0]  dataBusIn,
                output [7:0] dataBusOut,
    input RD,
    input WR,
    input sClk, 
    input [7:0] entera,   
    input [7:0] enterd,
    input clk2
    
    );
    
    reg [7:0] blockMem [255:0];
    //reg [7:0]outHold;
    
               //assign DataBus  = (RD)?blockMem[Address] : 8'hzz;
    assign dataBusOut = blockMem[Address]; 
    
 /*   always @(posedge clk2)
    begin
        blockMem[entera] <= enterd;
    end */
    
/*    always @(posedge sClk )begin
        if (WR) 
            //blockMem[Address] <= DataBus;
            blockMem[Address] <= dataBusIn;
    end */
    
    always @(*)
    begin
    if(sClk)
    begin
        if (WR) 
            blockMem[Address] <= dataBusIn;
    end 
    else if(clk2)
    begin
        blockMem[entera] <= enterd;
    end    
               
    end 
        
    
   /* initial begin
        //$readmemb("C:/Users/prasanna/Desktop/latest/Behavioural_YES_FPGA_No.srcs/sim_1/imports/Desktop/output.txt",blockMem);
            //$readmemb("/home/abhimanyu/Desktop/BiswasProject/latest/Behavioural_YES_FPGA_No.srcs/sim_1/imports/Desktop/output.txt",blockMem);
        
        blockMem[0] =  8'h00;
        blockMem[1] =  8'h00;
        blockMem[2] =  8'h00;
        blockMem[3] =  8'h00;
        blockMem[4] =  8'h00;
        blockMem[5] =  8'h00;
        blockMem[6] =  8'h00;
        blockMem[7] =  8'h00;
        blockMem[8] =  8'h00;
        blockMem[9] =  8'h00;
        blockMem[10] = 8'h00;
        blockMem[11] = 8'h00;
        blockMem[12] = 8'h00;
        blockMem[13] = 8'h00;
        blockMem[14] = 8'h00;
        blockMem[15] = 8'h00;
        blockMem[16] = 8'h00;
        blockMem[17] = 8'h00;
        blockMem[18] = 8'h00;
        blockMem[19] = 8'h00;
        blockMem[20] = 8'h00;
        blockMem[21] = 8'h00;
        blockMem[22] = 8'h00;
        blockMem[23] = 8'h00;
        blockMem[24] = 8'h00;
        blockMem[25] = 8'h00;
        blockMem[26] = 8'h0;
        blockMem[27] = 8'h0;
        blockMem[28] = 8'h0;
        blockMem[29] = 8'h0;
        blockMem[30] = 8'h0;
        blockMem[31] = 8'h0;
        blockMem[32] = 8'h0;
        blockMem[33] = 8'h0;
        blockMem[34] = 8'h0;
        blockMem[35] = 8'h0;
        blockMem[36] = 8'h0;
        blockMem[37] = 8'h0;
        blockMem[38] = 8'h0;
        blockMem[39] = 8'h0;
        blockMem[40] = 8'h0;
        blockMem[41] = 8'h0;
        blockMem[42] = 8'h0;
        blockMem[43] = 8'h0;
        blockMem[44] = 8'h0;
        blockMem[45] = 8'h0;
        blockMem[46] = 8'h0;
        blockMem[47] = 8'h0;
        blockMem[48] = 8'h0;
        blockMem[49] = 8'h0;
        blockMem[50] = 8'h0;
        blockMem[51] = 8'h0;
        blockMem[52] = 8'h0;
        blockMem[53] = 8'h0;
        blockMem[54] = 8'h0;
        blockMem[55] = 8'h0;
        blockMem[56] = 8'h0;
        blockMem[57] = 8'h0;
        blockMem[58] = 8'h0;
        blockMem[59] = 8'h0;
        blockMem[60] = 8'h0;
        blockMem[61] = 8'h0;
        blockMem[62] = 8'h0;
        blockMem[63] = 8'h0;
        blockMem[64] = 8'h0;
        blockMem[65] = 8'h0;
        blockMem[66] = 8'h0;
        blockMem[67] = 8'h0;
        blockMem[68] = 8'h0;
        blockMem[69] = 8'h0;
        blockMem[70] = 8'h0;
        blockMem[71] = 8'h0;
        blockMem[72] = 8'h0;
        blockMem[73] = 8'h0;
        blockMem[74] = 8'h0;
        blockMem[75] = 8'h0;
        blockMem[76] = 8'h0;
        blockMem[77] = 8'h0;
        blockMem[78] = 8'h0;
        blockMem[79] = 8'h0;
        blockMem[80] = 8'h0;
        blockMem[81] = 8'h0;
        blockMem[82] = 8'h0;
        blockMem[83] = 8'h0;
        blockMem[84] = 8'h0;
        blockMem[85] = 8'h0;
        blockMem[86] = 8'h0;
        blockMem[87] = 8'h0;
        blockMem[88] = 8'h0;
        blockMem[89] = 8'h0;
        blockMem[90] = 8'h0;
        blockMem[91] = 8'h0;
        blockMem[92] = 8'h0;
        blockMem[93] = 8'h0;
        blockMem[94] = 8'h0;
        blockMem[95] = 8'h0;
        blockMem[96] = 8'h0;
        blockMem[97] = 8'h0;
        blockMem[98] = 8'h0;
        blockMem[99] = 8'h0;
        blockMem[100] =8'h0;
        blockMem[101] =8'h0;
        blockMem[102] =8'h0;
        blockMem[103] =8'h0;
        blockMem[104] =8'h0;
        blockMem[105] =8'h0;
        blockMem[106] =8'h0;
        blockMem[107] =8'h0;
        blockMem[108] =8'h0;
        blockMem[109] =8'h0;
        blockMem[110] =8'h0;
        blockMem[111] =8'h0;
        blockMem[112] =8'h0;
        blockMem[113] =8'h0;
        blockMem[114] =8'h0;
        blockMem[115] =8'h0;
        blockMem[116] =8'h0;
        blockMem[117] =8'h0;
        blockMem[118] =8'h0;
        blockMem[119] =8'h0;
        blockMem[120] =8'h0;
        blockMem[121] =8'h0;
        blockMem[122] =8'h0;
        blockMem[123] =8'h0;
        blockMem[124] =8'h0;
        blockMem[125] =8'h0;
        blockMem[126] =8'h0;
        blockMem[127] =8'h0;
        blockMem[128] =8'h0;
        blockMem[129] =8'h0;
        blockMem[130] =8'h0;
        blockMem[131] =8'h0;
        blockMem[132] =8'h0;
        blockMem[133] =8'h0;
        blockMem[134] =8'h0;
        blockMem[135] =8'h0;
        blockMem[136] =8'h0;
        blockMem[137] =8'h0;
        blockMem[138] =8'h0;
        blockMem[139] =8'h0;
        blockMem[140] =8'h0;
        blockMem[141] =8'h0;
        blockMem[142] =8'h0;
        blockMem[143] =8'h0;
        blockMem[144] =8'h0;
        blockMem[145] =8'h0;
        blockMem[146] =8'h0;
        blockMem[147] =8'h0;
        blockMem[148] =8'h0;
        blockMem[149] =8'h0;
        blockMem[150] =8'h0;
        blockMem[151] =8'h0;
        blockMem[152] =8'h0;
        blockMem[153] =8'h0;
        blockMem[154] =8'h0;
        blockMem[155] =8'h0;
        blockMem[156] =8'h0;
        blockMem[157] =8'h0;
        blockMem[158] =8'h0;
        blockMem[159] =8'h0;
        blockMem[160] =8'h0;
        blockMem[161] =8'h0;
        blockMem[162] =8'h0;
        blockMem[163] =8'h0;
        blockMem[164] =8'h0;
        blockMem[165] =8'h0;
        blockMem[166] =8'h0;
        blockMem[167] =8'h0;
        blockMem[168] =8'h0;
        blockMem[169] =8'h0;
        blockMem[170] =8'h0;
        blockMem[171] =8'h0;
        blockMem[172] =8'h0;
        blockMem[173] =8'h0;
        blockMem[174] =8'h0;
        blockMem[175] =8'h0;
        blockMem[176] =8'h0;
        blockMem[177] =8'h0;
        blockMem[178] =8'h0;
        blockMem[179] =8'h0;
        blockMem[180] =8'h0;
        blockMem[181] =8'h0;
        blockMem[182] =8'h0;
        blockMem[183] =8'h0;
        blockMem[184] =8'h0;
        blockMem[185] =8'h0;
        blockMem[186] =8'h0;
        blockMem[187] =8'h0;
        blockMem[188] =8'h0;
        blockMem[189] =8'h0;
        blockMem[190] =8'h0;
        blockMem[191] =8'h0;
        blockMem[192] =8'h0;
        blockMem[193] =8'h0;
        blockMem[194] =8'h0;
        blockMem[195] =8'h0;
        blockMem[196] =8'h0;
        blockMem[197] =8'h0;
        blockMem[198] =8'h0;
        blockMem[199] =8'h0;
        blockMem[200] =8'h0;
        blockMem[201] =8'h0;
        blockMem[202] =8'h0;
        blockMem[203] =8'h0;
        blockMem[204] =8'h0;
        blockMem[205] =8'h0;
        blockMem[206] =8'h0;
        blockMem[207] =8'h0;
        blockMem[208] =8'h0;
        blockMem[209] =8'h0;
        blockMem[210] =8'h0;
        blockMem[211] =8'h0;
        blockMem[212] =8'h0;
        blockMem[213] =8'h0;
        blockMem[214] =8'h0;
        blockMem[215] =8'h0;
        blockMem[216] =8'h0;
        blockMem[217] =8'h0;
        blockMem[218] =8'h0;
        blockMem[219] =8'h0;
        blockMem[220] =8'h0;
        blockMem[221] =8'h0;
        blockMem[222] =8'h0;
        blockMem[223] =8'h0;
        blockMem[224] =8'h0;
        blockMem[225] =8'h0;
        blockMem[226] =8'h0;
        blockMem[227] =8'h0;
        blockMem[228] =8'h0;
        blockMem[229] =8'h0;
        blockMem[230] =8'h0;
        blockMem[231] =8'h0;
        blockMem[232] =8'h0;
        blockMem[233] =8'h0;
        blockMem[234] =8'h0;
        blockMem[235] =8'h0;
        blockMem[236] =8'h0;
        blockMem[237] =8'h0;
        blockMem[238] =8'h0;
        blockMem[239] =8'h0;
        blockMem[240] =8'h0;
        blockMem[241] =8'h0;
        blockMem[242] =8'h0;
        blockMem[243] =8'h0;
        blockMem[244] =8'h0;
        blockMem[245] =8'h0;
        blockMem[246] =8'h0;
        blockMem[247] =8'h0;
        blockMem[248] =8'h0;
        blockMem[249] =8'h0;
        blockMem[250] =8'h0;
        blockMem[251] =8'h0;
        blockMem[252] =8'h0;
        blockMem[253] =8'h0;
        blockMem[254] =8'h0;
        blockMem[255] =8'h0; 
        
       
   // blockMem[0] = 8'h01;  //CLR
                blockMem[1] = 8'h1f;  //MVS<rn>
                blockMem[2] = 8'h62;  //STA<rn>
                blockMem[3] = 8'h9c;  //SBI<rn><od>
                blockMem[4] = 8'h54;  //DCR<rn>
                blockMem[5] = 8'he5;  //XRA<rn>
                blockMem[6] = 8'hb2;  //SCA<rn>
                blockMem[7] = 8'h62;  //STA<rn>
                blockMem[8] = 8'hb6;  //SCA<rn>
                blockMem[9] = 8'h47;  //INC<rn>
                blockMem[10] = 8'h58;  //MVI<rn><od>
                blockMem[11] = 8'h5b;  //MVI<rn><od>
                blockMem[12] = 8'he4;  //XRA<rn>
                blockMem[13] = 8'hb6;  //SCA<rn>
                blockMem[14] = 8'h7d;  //POP<rn>
                blockMem[15] = 8'h7b;  //POP<rn>
                blockMem[16] = 8'h61;  //STA<rn>
                blockMem[17] = 8'h79;  //POP<rn>
                blockMem[18] = 8'h5e;  //MVI<rn><od>
                blockMem[19] = 8'h13;  //MVD<rn>
                blockMem[20] = 8'h86;  //ADA<rn>
                blockMem[21] = 8'h83;  //ADA<rn>
                blockMem[22] = 8'h58;  //MVI<rn><od>
                blockMem[23] = 8'hed;  //XRI<rn><od>
                blockMem[24] = 8'h6f;  //PSH<rn>
                blockMem[25] = 8'hcc;  //ANI<rn><od>
                blockMem[26] = 8'h18;  //RSP
                blockMem[27] = 8'hea;  //XRI<rn><od>
                blockMem[28] = 8'h5a;  //MVI<rn><od>
                blockMem[29] = 8'h59;  //MVI<rn><od>
                blockMem[30] = 8'h1f;  //MVS<rn>
                blockMem[31] = 8'h00;  //SBA<rn>
                blockMem[32] = 8'hdd;  //ORI<rn><od>
                blockMem[33] = 8'h22;  //NOT<rn>
                blockMem[34] = 8'h6c;  //PSH<rn>
                blockMem[35] = 8'h6d;  //PSH<rn>
                blockMem[36] = 8'h62;  //STA<rn>
                blockMem[37] = 8'h5e;  //MVI<rn><od>
                blockMem[38] = 8'h8d;  //ADI<rn><od>
                blockMem[39] = 8'h9b;  //SBI<rn><od>
                blockMem[40] = 8'h11;  //MVD<rn>
                blockMem[41] = 8'h00;  //ACA<rn>
                blockMem[42] = 8'h76;  //LDA<rn>
                blockMem[43] = 8'he6;  //XRA<rn>
                blockMem[44] = 8'h77;  //LDA<rn>
                blockMem[45] = 8'h71;  //LDA<rn>
                blockMem[46] = 8'hd9;  //ORI<rn><od>
                blockMem[47] = 8'h17;  //MVD<rn>
                blockMem[48] = 8'h67;  //STA<rn>
                blockMem[49] = 8'h97;  //SBA<rn>
                blockMem[50] = 8'h24;  //NOT<rn>
                blockMem[51] = 8'h19;  //MVS<rn>
                blockMem[52] = 8'h71;  //LDA<rn>
                blockMem[53] = 8'h61;  //STA<rn>
                blockMem[54] = 8'h6c;  //PSH<rn>
                blockMem[55] = 8'h61;  //STA<rn>
                blockMem[56] = 8'h1a;  //MVS<rn>
                blockMem[57] = 8'ha3;  //ACA<rn>
                blockMem[58] = 8'hdb;  //ORI<rn><od>
                blockMem[59] = 8'h13;  //MVD<rn>
                blockMem[60] = 8'h58;  //MVI<rn><od>
                blockMem[61] = 8'h68;  //PSH<rn>
                blockMem[62] = 8'h14;  //MVD<rn>
                blockMem[63] = 8'hbe;  //SCI<rn><od>
                blockMem[64] = 8'hc8;  //ANI<rn><od>
                blockMem[65] = 8'h6a;  //PSH<rn>
                blockMem[66] = 8'h57;  //DCR<rn>
                blockMem[67] = 8'h22;  //NOT<rn>
                blockMem[68] = 8'h67;  //STA<rn>
                blockMem[69] = 8'haf;  //ACI<rn><od>
                blockMem[70] = 8'h5c;  //MVI<rn><od>
                blockMem[71] = 8'h5d;  //MVI<rn><od>
                blockMem[72] = 8'h6f;  //PSH<rn>
                blockMem[73] = 8'h6c;  //PSH<rn>
                blockMem[74] = 8'hbb;  //SCI<rn><od>
                blockMem[75] = 8'h7d;  //POP<rn>
                blockMem[76] = 8'hd8;  //ORI<rn><od>
                blockMem[77] = 8'h68;  //PSH<rn>
                blockMem[78] = 8'h7c;  //POP<rn>
                blockMem[79] = 8'h77;  //LDA<rn>
                blockMem[80] = 8'h58;  //MVI<rn><od>
                blockMem[81] = 8'h7f;  //POP<rn>
                blockMem[82] = 8'h13;  //MVD<rn>
                blockMem[83] = 8'hde;  //ORI<rn><od>
                blockMem[84] = 8'h71;  //LDA<rn>
                blockMem[85] = 8'h8e;  //ADI<rn><od>
                blockMem[86] = 8'h42;  //INC<rn>
                blockMem[87] = 8'h6a;  //PSH<rn>
                blockMem[88] = 8'ha5;  //ACA<rn>
                blockMem[89] = 8'hd6;  //ORA<rn>
                blockMem[90] = 8'h11;  //MVD<rn>
                blockMem[91] = 8'h63;  //STA<rn>
                blockMem[92] = 8'hd2;  //ORA<rn>
                blockMem[93] = 8'hc3;  //ANA<rn>
                blockMem[94] = 8'h11;  //MVD<rn>
                blockMem[95] = 8'h62;  //STA<rn>
                blockMem[96] = 8'hb4;  //SCA<rn>
                blockMem[97] = 8'h66;  //STA<rn>
                blockMem[98] = 8'hd0;  //ORA<rn>
                blockMem[99] = 8'h6a;  //PSH<rn>
                blockMem[100] = 8'h69;  //PSH<rn>
                blockMem[101] = 8'h1d;  //MVS<rn>
                blockMem[102] = 8'ha2;  //ACA<rn>
                blockMem[103] = 8'heb;  //XRI<rn><od>
                blockMem[104] = 8'h54;  //DCR<rn>
                blockMem[105] = 8'h19;  //MVS<rn>
                blockMem[106] = 8'h5a;  //MVI<rn><od>
                blockMem[107] = 8'hbc;  //SCI<rn><od>
                blockMem[108] = 8'h93;  //SBA<rn>
                blockMem[109] = 8'he8;  //XRI<rn><od>
                blockMem[110] = 8'h69;  //PSH<rn>
                blockMem[111] = 8'h99;  //SBI<rn><od>
                blockMem[112] = 8'h7d;  //POP<rn>
                blockMem[113] = 8'ha7;  //ACA<rn>
                blockMem[114] = 8'h26;  //NOT<rn>
                blockMem[115] = 8'h91;  //SBA<rn>
                blockMem[116] = 8'hbe;  //SCI<rn><od>
                blockMem[117] = 8'h6a;  //PSH<rn>
                blockMem[118] = 8'hd5;  //ORA<rn>
                blockMem[119] = 8'hc4;  //ANA<rn>
                blockMem[120] = 8'h66;  //STA<rn>
                blockMem[121] = 8'h79;  //POP<rn>
                blockMem[122] = 8'h61;  //STA<rn>
                blockMem[123] = 8'hb2;  //SCA<rn>
                blockMem[124] = 8'hc3;  //ANA<rn>
                blockMem[125] = 8'h7e;  //POP<rn>
                blockMem[126] = 8'h6d;  //PSH<rn>
                blockMem[127] = 8'h97;  //SBA<rn>
                blockMem[128] = 8'h6f;  //PSH<rn>
                blockMem[129] = 8'haa;  //ACI<rn><od>
                blockMem[130] = 8'h00;  //ACA<rn>
                blockMem[131] = 8'h61;  //STA<rn>
                blockMem[132] = 8'h96;  //SBA<rn>
                blockMem[133] = 8'he9;  //XRI<rn><od>
                blockMem[134] = 8'h65;  //STA<rn>
                blockMem[135] = 8'h61;  //STA<rn>
                blockMem[136] = 8'h10;  //LSP
                blockMem[137] = 8'h7d;  //POP<rn>
                blockMem[138] = 8'h17;  //MVD<rn>
                blockMem[139] = 8'h58;  //MVI<rn><od>
                blockMem[140] = 8'h66;  //STA<rn>
                blockMem[141] = 8'h7a;  //POP<rn>
                blockMem[142] = 8'h79;  //POP<rn>
                blockMem[143] = 8'h7b;  //POP<rn>
                blockMem[144] = 8'h11;  //MVD<rn>
                blockMem[145] = 8'h69;  //PSH<rn>
                blockMem[146] = 8'hd3;  //ORA<rn>
                blockMem[147] = 8'h7f;  //POP<rn>
                blockMem[148] = 8'h20;  //NOT<rn>
                blockMem[149] = 8'h6a;  //PSH<rn>
                blockMem[150] = 8'h7a;  //POP<rn>
                blockMem[151] = 8'h5c;  //MVI<rn><od>
                blockMem[152] = 8'h27;  //NOT<rn>
                blockMem[153] = 8'h1c;  //MVS<rn>
                blockMem[154] = 8'h6f;  //PSH<rn>
                blockMem[155] = 8'h61;  //STA<rn>
                blockMem[156] = 8'hc3;  //ANA<rn>
                blockMem[157] = 8'hef;  //XRI<rn><od>
                blockMem[158] = 8'h68;  //PSH<rn>
                blockMem[159] = 8'h78;  //POP<rn>
                blockMem[160] = 8'h40;  //INC<rn>
                blockMem[161] = 8'h98;  //SBI<rn><od>
                blockMem[162] = 8'h6a;  //PSH<rn>
                blockMem[163] = 8'h7d;  //POP<rn>
                blockMem[164] = 8'h65;  //STA<rn>
                blockMem[165] = 8'h1d;  //MVS<rn>
                blockMem[166] = 8'hbf;  //SCI<rn><od>
                blockMem[167] = 8'h6b;  //PSH<rn>
                blockMem[168] = 8'h73;  //LDA<rn>
                blockMem[169] = 8'h55;  //DCR<rn>
                blockMem[170] = 8'hbb;  //SCI<rn><od>
                blockMem[171] = 8'hc2;  //ANA<rn>
                blockMem[172] = 8'h73;  //LDA<rn>
                blockMem[173] = 8'hd3;  //ORA<rn>
                blockMem[174] = 8'h58;  //MVI<rn><od>
                blockMem[175] = 8'h67;  //STA<rn>
                blockMem[176] = 8'h5d;  //MVI<rn><od>
                blockMem[177] = 8'h25;  //NOT<rn>
                blockMem[178] = 8'h5e;  //MVI<rn><od>
                blockMem[179] = 8'h40;  //INC<rn>
                blockMem[180] = 8'h7c;  //POP<rn>
                blockMem[181] = 8'h1f;  //MVS<rn>
                blockMem[182] = 8'h6e;  //PSH<rn>
                blockMem[183] = 8'hdf;  //ORI<rn><od>
                blockMem[184] = 8'hce;  //ANI<rn><od>
                blockMem[185] = 8'h63;  //STA<rn>
                blockMem[186] = 8'h5d;  //MVI<rn><od>
                blockMem[187] = 8'hcc;  //ANI<rn><od>
                blockMem[188] = 8'h5d;  //MVI<rn><od>
                blockMem[189] = 8'h43;  //INC<rn>
                blockMem[190] = 8'h51;  //DCR<rn>
                blockMem[191] = 8'h76;  //LDA<rn>
                blockMem[192] = 8'h6f;  //PSH<rn>
                blockMem[193] = 8'h14;  //MVD<rn>
                blockMem[194] = 8'h59;  //MVI<rn><od>
                blockMem[195] = 8'h62;  //STA<rn>
                blockMem[196] = 8'hde;  //ORI<rn><od>
                blockMem[197] = 8'h51;  //DCR<rn>
                blockMem[198] = 8'h5e;  //MVI<rn><od>
                blockMem[199] = 8'h6a;  //PSH<rn>
                blockMem[200] = 8'h62;  //STA<rn>
                blockMem[201] = 8'h73;  //LDA<rn>
                blockMem[202] = 8'h69;  //PSH<rn>
                blockMem[203] = 8'h7a;  //POP<rn>
                blockMem[204] = 8'h64;  //STA<rn>
                blockMem[205] = 8'h76;  //LDA<rn>
                blockMem[206] = 8'h1b;  //MVS<rn>
                blockMem[207] = 8'h58;  //MVI<rn><od>
                blockMem[208] = 8'h69;  //PSH<rn>
                blockMem[209] = 8'h78;  //POP<rn>
                blockMem[210] = 8'h1a;  //MVS<rn>
                blockMem[211] = 8'h9e;  //SBI<rn><od>
                blockMem[212] = 8'h94;  //SBA<rn>
                blockMem[213] = 8'h78;  //POP<rn>
                blockMem[214] = 8'h92;  //SBA<rn>
                blockMem[215] = 8'h65;  //STA<rn>
                blockMem[216] = 8'h20;  //NOT<rn>
                blockMem[217] = 8'h7a;  //POP<rn>
                blockMem[218] = 8'h77;  //LDA<rn>
                blockMem[219] = 8'h2;  //CLC
                blockMem[220] = 8'h59;  //MVI<rn><od>
                blockMem[221] = 8'h77;  //LDA<rn>
                blockMem[222] = 8'h5b;  //MVI<rn><od>
                blockMem[223] = 8'h00;  //ACA<rn>
                blockMem[224] = 8'h66;  //STA<rn>
                blockMem[225] = 8'h8a;  //ADI<rn><od>
                blockMem[226] = 8'h17;  //MVD<rn>
                blockMem[227] = 8'hec;  //XRI<rn><od>
                blockMem[228] = 8'h5d;  //MVI<rn><od>
                blockMem[229] = 8'h59;  //MVI<rn><od>
                blockMem[230] = 8'he7;  //XRA<rn>
                blockMem[231] = 8'h1a;  //MVS<rn>
                blockMem[232] = 8'h74;  //LDA<rn>
                blockMem[233] = 8'h5d;  //MVI<rn><od>
                blockMem[234] = 8'h88;  //ADI<rn><od>
                blockMem[235] = 8'h1b;  //MVS<rn>
                blockMem[236] = 8'h15;  //MVD<rn>
                blockMem[237] = 8'h67;  //STA<rn>
                blockMem[238] = 8'h77;  //LDA<rn>
                blockMem[239] = 8'h42;  //INC<rn>
                blockMem[240] = 8'he1;  //XRA<rn>
                blockMem[241] = 8'h66;  //STA<rn>
                blockMem[242] = 8'hbe;  //SCI<rn><od>
                blockMem[243] = 8'h41;  //INC<rn>
                blockMem[244] = 8'hce;  //ANI<rn><od>
                blockMem[245] = 8'h45;  //INC<rn>
                blockMem[246] = 8'h7f;  //POP<rn>
                blockMem[247] = 8'h88;  //ADI<rn><od>
                blockMem[248] = 8'h53;  //DCR<rn>
                blockMem[249] = 8'h79;  //POP<rn>
                blockMem[250] = 8'h6d;  //PSH<rn>
                blockMem[251] = 8'h62;  //STA<rn>
                blockMem[252] = 8'h9a;  //SBI<rn><od>
                blockMem[253] = 8'hef;  //XRI<rn><od>
                blockMem[254] = 8'h7c;  //POP<rn>
                blockMem[255] = 8'h01; //CLR
*/

 //   end 
    
endmodule